library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- This file simulates a 512x8 synchronous RAM component.
-- The program to be executed is encoded by initializing the "mem_data" signal (see below).

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_arith.all;
USE IEEE.std_logic_unsigned.all;

entity microram_sim is
port (  CLOCK   : in STD_LOGIC ;
		ADDRESS	: in STD_LOGIC_VECTOR (8 downto 0);
		DATAOUT : out STD_LOGIC_VECTOR (7 downto 0);
		DATAIN  : in STD_LOGIC_VECTOR (7 downto 0);
		WE	: in STD_LOGIC 
	);
end entity microram_sim;

architecture a of microram_sim is
type t_mem_data is array(0 to 511) of std_logic_vector(7 downto 0);

-- Your program is entered here, as initialization values for the "mem_data" signal.
signal mem_data : t_mem_data := (0 => "11110000", -- CLR A (dummy first instruction)
                                 1 => "00000000", -- LOAD 10,A  
                                 2 => X"0A",      -- ADDRESS -> 10
	                             3 => "00010000", -- BCDO A       
	                             4 => "10100000", -- LSL A       
	                             5 => "00010000", -- BCDO A 
	                             6 => "00000001", -- LOAD 11,B  
	                             7 => X"0B",      -- ADDRESS -> 11
	                           	 8 => "10000000", -- ADD A 
	                           	 9 => "00010000", -- BCDO A       
	                    	     -- test data --
                                10 => "00000001", -- memory location 10 set to 1
                                11 => "00000101", -- memory location 11 set to 5
                            others => "11110000"); -- all other memory locations set to CLR A instr

--signal mem_data : t_mem_data := (0 => "11110000", -- CLR A (dummy first instruction)
--                                 1 => "00000000", -- LOAD 10,A  
--                                 2 => X"0A",      -- ADDRESS -> 10
--	                             3 => "00001000", -- OUT A       
--	                             4 => "10100000", -- LSL A       
--	                             5 => "00001000", -- OUT A 
--	                             6 => "00000001", -- LOAD 11,B  
--	                             7 => X"0B",      -- ADDRESS -> 11
--	                           	 8 => "10000000", -- ADD A 
--	                           	 9 => "00001000", -- OUT A       
--	                    	     -- test data --
--                                10 => "00000001", -- memory location 10 set to 1
--                                11 => "00000101", -- memory location 11 set to 5
--                            others => "11110000"); -- all other memory locations set to CLR A instr

begin
RAM_Process : process(CLOCK)
variable memaddr : INTEGER range 0 to 511;
begin
  if(rising_edge(CLOCK)) then
     memaddr := CONV_INTEGER(ADDRESS);
     if(we='1') then
        mem_data(memaddr) <= DATAIN;
        DATAOUT <= DATAIN;
     else
        DATAOUT <= mem_data(memaddr);
     end if;
  end if;
end process;
end architecture a;

